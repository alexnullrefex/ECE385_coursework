module Multiplier();



endmodule